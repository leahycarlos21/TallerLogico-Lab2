module and_(input a, input b,
				output c);

//Implica logica combinacional
assign c = a & b;
				
endmodule

// a| b, !a