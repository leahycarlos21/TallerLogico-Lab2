module not_(input a, output b);
assign b = !a;
endmodule
