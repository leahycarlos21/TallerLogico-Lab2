module xor_(input a, input b,
				output c);

//assign c = a ^ b;
//assign c = (!a & b) | (a & !b);

//empieza

//logic w;
//
//always_comb begin
//	w = a ^ b;
//end
//
//assign c = w;

//termina


logic w1, w2, w3, w4;

not_ N1(a,w1);
not_ N2(b, w2);

and_ A1(b, w1, w3);
and_ A2(w2, a, w4);

or_ O1(w3, w4, c);
 
endmodule
