ENTITY adder4bit IS 
PORT (a0: IN BIT;	--Primer numero
		a1: IN BIT;
		a2: IN BIT;
		a3: IN BIT;
		b0: IN BIT;	--Segundo numero
		b1: IN BIT;
		b2: IN BIT;
		b3: IN BIT;
		c0: IN BIT;	--acarreo inicail
		s0: OUT BIT;--Resultado
		s1: OUT BIT;
		s2: OUT BIT;
		s3: OUT BIT;
		cout: OUT BIT
		);
END ENTITY adder4bit;

ARCHITECTURE adder4bit_arch OF adder4bit IS

COMPONENT fulladder_ent
	PORT (a: IN BIT;
			b: IN BIT;		
			cin: IN BIT;
			sum: OUT BIT;
			cout: OUT BIT
			);
END COMPONENT;

SIGNAL c1, c2, c3: BIT:= '0';
BEGIN
	fa0: fulladder_ent port map(
										a => a0,
										b => b0,
										cin => c0,
										sum => s0,
										cout => c1);
	fa1: fulladder_ent port map(
										a => a1,
										b => b1,
										cin => c1,
										sum => s1,
										cout => c2
										);
	fa2: fulladder_ent port map(
										a => a2,
										b => b2,
										cin => c2,
										sum => s2,
										cout => c3
										);
	fa3: fulladder_ent port map(
										a => a3,
										b => b3,
										cin => c3,
										sum => s3,
										cout => cout
										);
										
END ARCHITECTURE adder4bit_arch;